
class top_sqr extends uvm_sequencer;
  `uvm_component_utils(top_sqr)
  `new_component
  
  apb_sqr sqr_inst;
endclass