typedef uvm_sequencer#(axi_tx) axi_sqr;


