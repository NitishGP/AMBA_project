
class axi_tx extends uvm_sequence_item;
	`NEW_OBJ

	`uvm_object_utils_begin(axi_tx)
	`uvm_object_utils_end
endclass
