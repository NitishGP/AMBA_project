
class axi_base_seq extends uvm_sequence#(axi_tx);
	`uvm_object_utils(axi_base_seq)
	`NEW_OBJ

	task pre_body();
	endtask

	task post_body();
	endtask
endclass


