class axi_res extends uvm_component;
	`uvm_component_utils(axi_res)
	`NEW_COMP
	
	function void build();
	endfunction

	task run();
	endtask
endclass
