
interface axi_intf(input reg clk,rst);
	
endinterface
